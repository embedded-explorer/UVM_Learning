//--------------------------------------------------------------------
// UVM Transaction Example
// Package
//--------------------------------------------------------------------

package my_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  `include "my_sequence_item.sv"
  `include "my_test.sv"

endpackage
